

module  tb_memory_rw();


wire    a;
wire    b;

reg     x;
reg     y;

initial begin
    
//  LEER ARCHIVO DE SEÑAL Y MANDARLO A LA MEMORIA RAM

//  PRUEBAS DE ESTADOS DE AUTOMATA

//  EMISION DE SEÑAL CAPTURADA


end


endmodule
